`include "uart_if.sv"
module rx_checker_module (uart_io uart);

    

    
    // property check_rx_done_prop;
    //   @(posedge uart.clk)
    // endproperty

    // AP_RX_DONE : assert property (check_rx_done_prop);  
endmodule