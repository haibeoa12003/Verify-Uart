`define FREQUENCY 50000000
`define BAURATE 115200